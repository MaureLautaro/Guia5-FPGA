// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
// Created on Mon Nov 03 21:46:32 2025

// synthesis message_off 10175

`timescale 1ns/1ns

module I2C (
    reset,clock,SDA,fin_dir,fin_dato,soy);

    input reset;
    input clock;
    input SDA;
    input fin_dir;
    input fin_dato;
    input soy;
    tri0 reset;
    tri0 SDA;
    tri0 fin_dir;
    tri0 fin_dato;
    tri0 soy;
    reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter ocioso=0,RW=1,Guardardir=2,GuardarDato=3,ACK=4;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or SDA or fin_dir or fin_dato or soy)
    begin
        if (reset) begin
            reg_fstate <= ocioso;
        end
        else begin
            case (fstate)
                ocioso: begin
                    if ((SDA == 1'b0))
                        reg_fstate <= Guardardir;
                    else if ((SDA == 1'b1))
                        reg_fstate <= ocioso;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= ocioso;
                end
                RW: begin
                    reg_fstate <= ACK;
                end
                Guardardir: begin
                    if (((fin_dir == 1'b1) | (soy == 1'b0)))
                        reg_fstate <= ocioso;
                    else if (((fin_dir == 1'b1) | (soy == 1'b1)))
                        reg_fstate <= RW;
                    else if ((fin_dir == 1'b0))
                        reg_fstate <= Guardardir;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= Guardardir;
                end
                GuardarDato: begin
                    if ((fin_dato == 1'b0))
                        reg_fstate <= GuardarDato;
                    else if ((fin_dato == 1'b1))
                        reg_fstate <= ocioso;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= GuardarDato;
                end
                ACK: begin
                    reg_fstate <= GuardarDato;
                end
                default: begin
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // I2C

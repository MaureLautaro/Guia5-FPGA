-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Oct 30 20:59:26 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY I2C IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        SDA : IN STD_LOGIC := '0';
        fin_dir : IN STD_LOGIC := '0';
        fin_dato : IN STD_LOGIC := '0';
        soy : IN STD_LOGIC := '0'
    );
END I2C;

ARCHITECTURE BEHAVIOR OF I2C IS
    TYPE type_fstate IS (ocioso,RW,Guardardir,GuardarDato,ACK);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,SDA,fin_dir,fin_dato,soy)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= ocioso;
        ELSE
            CASE fstate IS
                WHEN ocioso =>
                    IF ((SDA = '0')) THEN
                        reg_fstate <= Guardardir;
                    ELSIF ((SDA = '1')) THEN
                        reg_fstate <= ocioso;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ocioso;
                    END IF;
                WHEN RW =>
                    reg_fstate <= ACK;
                WHEN Guardardir =>
                    IF (((fin_dir = '1') OR (soy = '0'))) THEN
                        reg_fstate <= ocioso;
                    ELSIF (((fin_dir = '1') OR (soy = '1'))) THEN
                        reg_fstate <= RW;
                    ELSIF ((fin_dir = '0')) THEN
                        reg_fstate <= Guardardir;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guardardir;
                    END IF;
                WHEN GuardarDato =>
                    IF ((fin_dato = '0')) THEN
                        reg_fstate <= GuardarDato;
                    ELSIF ((fin_dato = '1')) THEN
                        reg_fstate <= ocioso;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= GuardarDato;
                    END IF;
                WHEN ACK =>
                    reg_fstate <= GuardarDato;
                WHEN OTHERS => 
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;

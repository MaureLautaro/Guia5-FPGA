-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Wed Oct 29 20:27:44 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY mult2x2_Ca2 IS 
	PORT
	(
		A1 :  IN  STD_LOGIC;
		A0 :  IN  STD_LOGIC;
		B0 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		clk :  IN  STD_LOGIC;
		V :  OUT  STD_LOGIC;
		r0 :  OUT  STD_LOGIC;
		r1 :  OUT  STD_LOGIC;
		r2 :  OUT  STD_LOGIC;
		r3 :  OUT  STD_LOGIC
	);
END mult2x2_Ca2;

ARCHITECTURE bdf_type OF mult2x2_Ca2 IS 

COMPONENT sumador_completo
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 Cin : IN STD_LOGIC;
		 S : OUT STD_LOGIC;
		 Cout : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_40 <= '1';
SYNTHESIZED_WIRE_41 <= '1';
SYNTHESIZED_WIRE_24 <= '0';
SYNTHESIZED_WIRE_26 <= '1';
SYNTHESIZED_WIRE_27 <= '0';
SYNTHESIZED_WIRE_38 <= '0';



PROCESS(clk,SYNTHESIZED_WIRE_40,SYNTHESIZED_WIRE_40)
BEGIN
IF (SYNTHESIZED_WIRE_40 = '0') THEN
	SYNTHESIZED_WIRE_44 <= '0';
ELSIF (SYNTHESIZED_WIRE_40 = '0') THEN
	SYNTHESIZED_WIRE_44 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_44 <= A0;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_40,SYNTHESIZED_WIRE_40)
BEGIN
IF (SYNTHESIZED_WIRE_40 = '0') THEN
	SYNTHESIZED_WIRE_45 <= '0';
ELSIF (SYNTHESIZED_WIRE_40 = '0') THEN
	SYNTHESIZED_WIRE_45 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_45 <= A1;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_41,SYNTHESIZED_WIRE_41)
BEGIN
IF (SYNTHESIZED_WIRE_41 = '0') THEN
	r0 <= '0';
ELSIF (SYNTHESIZED_WIRE_41 = '0') THEN
	r0 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	r0 <= SYNTHESIZED_WIRE_5;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_41,SYNTHESIZED_WIRE_41)
BEGIN
IF (SYNTHESIZED_WIRE_41 = '0') THEN
	r1 <= '0';
ELSIF (SYNTHESIZED_WIRE_41 = '0') THEN
	r1 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	r1 <= SYNTHESIZED_WIRE_8;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_40,SYNTHESIZED_WIRE_40)
BEGIN
IF (SYNTHESIZED_WIRE_40 = '0') THEN
	SYNTHESIZED_WIRE_43 <= '0';
ELSIF (SYNTHESIZED_WIRE_40 = '0') THEN
	SYNTHESIZED_WIRE_43 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_43 <= B0;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_40,SYNTHESIZED_WIRE_40)
BEGIN
IF (SYNTHESIZED_WIRE_40 = '0') THEN
	SYNTHESIZED_WIRE_47 <= '0';
ELSIF (SYNTHESIZED_WIRE_40 = '0') THEN
	SYNTHESIZED_WIRE_47 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	SYNTHESIZED_WIRE_47 <= B1;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_41,SYNTHESIZED_WIRE_41)
BEGIN
IF (SYNTHESIZED_WIRE_41 = '0') THEN
	r2 <= '0';
ELSIF (SYNTHESIZED_WIRE_41 = '0') THEN
	r2 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	r2 <= SYNTHESIZED_WIRE_15;
END IF;
END PROCESS;


PROCESS(clk,SYNTHESIZED_WIRE_41,SYNTHESIZED_WIRE_41)
BEGIN
IF (SYNTHESIZED_WIRE_41 = '0') THEN
	r3 <= '0';
ELSIF (SYNTHESIZED_WIRE_41 = '0') THEN
	r3 <= '1';
ELSIF (RISING_EDGE(clk)) THEN
	r3 <= SYNTHESIZED_WIRE_18;
END IF;
END PROCESS;


V <= SYNTHESIZED_WIRE_42 XOR SYNTHESIZED_WIRE_21;


SYNTHESIZED_WIRE_5 <= SYNTHESIZED_WIRE_43 AND SYNTHESIZED_WIRE_44;


SYNTHESIZED_WIRE_48 <= NOT(SYNTHESIZED_WIRE_45);



SYNTHESIZED_WIRE_25 <= NOT(SYNTHESIZED_WIRE_44);



b2v_inst12 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_46,
		 B => SYNTHESIZED_WIRE_23,
		 Cin => SYNTHESIZED_WIRE_24,
		 S => SYNTHESIZED_WIRE_8,
		 Cout => SYNTHESIZED_WIRE_30);



b2v_inst14 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_25,
		 B => SYNTHESIZED_WIRE_26,
		 Cin => SYNTHESIZED_WIRE_27,
		 S => SYNTHESIZED_WIRE_35,
		 Cout => SYNTHESIZED_WIRE_39);



b2v_inst16 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_28,
		 B => SYNTHESIZED_WIRE_46,
		 Cin => SYNTHESIZED_WIRE_30,
		 S => SYNTHESIZED_WIRE_15,
		 Cout => SYNTHESIZED_WIRE_42);


b2v_inst17 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_31,
		 B => SYNTHESIZED_WIRE_46,
		 Cin => SYNTHESIZED_WIRE_42,
		 S => SYNTHESIZED_WIRE_18,
		 Cout => SYNTHESIZED_WIRE_21);



SYNTHESIZED_WIRE_46 <= SYNTHESIZED_WIRE_43 AND SYNTHESIZED_WIRE_45;


SYNTHESIZED_WIRE_28 <= SYNTHESIZED_WIRE_47 AND SYNTHESIZED_WIRE_34;


SYNTHESIZED_WIRE_23 <= SYNTHESIZED_WIRE_47 AND SYNTHESIZED_WIRE_35;


SYNTHESIZED_WIRE_31 <= SYNTHESIZED_WIRE_47 AND SYNTHESIZED_WIRE_48;


b2v_inst6 : sumador_completo
PORT MAP(A => SYNTHESIZED_WIRE_48,
		 B => SYNTHESIZED_WIRE_38,
		 Cin => SYNTHESIZED_WIRE_39,
		 S => SYNTHESIZED_WIRE_34);





END bdf_type;
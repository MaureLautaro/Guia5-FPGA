library verilog;
use verilog.vl_types.all;
entity mult2x2_vlg_vec_tst is
end mult2x2_vlg_vec_tst;
